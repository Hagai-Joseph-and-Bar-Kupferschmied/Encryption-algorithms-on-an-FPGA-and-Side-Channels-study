module sbox (
				input [7:0] originalByte, 
				output reg [7:0] subbedByte
			);


	always@(originalByte)
    begin
        case (originalByte)
         8'h00: subbedByte=8'h63;
		   8'h01: subbedByte=8'h7c;
		   8'h02: subbedByte=8'h77;
		   8'h03: subbedByte=8'h7b;
		   8'h04: subbedByte=8'hf2;
		   8'h05: subbedByte=8'h6b;
		   8'h06: subbedByte=8'h6f;
		   8'h07: subbedByte=8'hc5;
		   8'h08: subbedByte=8'h30;
		   8'h09: subbedByte=8'h01;
		   8'h0a: subbedByte=8'h67;
		   8'h0b: subbedByte=8'h2b;
		   8'h0c: subbedByte=8'hfe;
		   8'h0d: subbedByte=8'hd7;
		   8'h0e: subbedByte=8'hab;
		   8'h0f: subbedByte=8'h76;
		   8'h10: subbedByte=8'hca;
		   8'h11: subbedByte=8'h82;
		   8'h12: subbedByte=8'hc9;
		   8'h13: subbedByte=8'h7d;
		   8'h14: subbedByte=8'hfa;
		   8'h15: subbedByte=8'h59;
		   8'h16: subbedByte=8'h47;
		   8'h17: subbedByte=8'hf0;
		   8'h18: subbedByte=8'had;
		   8'h19: subbedByte=8'hd4;
		   8'h1a: subbedByte=8'ha2;
		   8'h1b: subbedByte=8'haf;
		   8'h1c: subbedByte=8'h9c;
		   8'h1d: subbedByte=8'ha4;
		   8'h1e: subbedByte=8'h72;
		   8'h1f: subbedByte=8'hc0;
		   8'h20: subbedByte=8'hb7;
		   8'h21: subbedByte=8'hfd;
		   8'h22: subbedByte=8'h93;
		   8'h23: subbedByte=8'h26;
		   8'h24: subbedByte=8'h36;
		   8'h25: subbedByte=8'h3f;
		   8'h26: subbedByte=8'hf7;
		   8'h27: subbedByte=8'hcc;
		   8'h28: subbedByte=8'h34;
		   8'h29: subbedByte=8'ha5;
		   8'h2a: subbedByte=8'he5;
		   8'h2b: subbedByte=8'hf1;
		   8'h2c: subbedByte=8'h71;
		   8'h2d: subbedByte=8'hd8;
		   8'h2e: subbedByte=8'h31;
		   8'h2f: subbedByte=8'h15;
		   8'h30: subbedByte=8'h04;
		   8'h31: subbedByte=8'hc7;
		   8'h32: subbedByte=8'h23;
		   8'h33: subbedByte=8'hc3;
		   8'h34: subbedByte=8'h18;
		   8'h35: subbedByte=8'h96;
		   8'h36: subbedByte=8'h05;
		   8'h37: subbedByte=8'h9a;
		   8'h38: subbedByte=8'h07;
		   8'h39: subbedByte=8'h12;
		   8'h3a: subbedByte=8'h80;
		   8'h3b: subbedByte=8'he2;
		   8'h3c: subbedByte=8'heb;
		   8'h3d: subbedByte=8'h27;
		   8'h3e: subbedByte=8'hb2;
		   8'h3f: subbedByte=8'h75;
		   8'h40: subbedByte=8'h09;
		   8'h41: subbedByte=8'h83;
		   8'h42: subbedByte=8'h2c;
		   8'h43: subbedByte=8'h1a;
		   8'h44: subbedByte=8'h1b;
		   8'h45: subbedByte=8'h6e;
		   8'h46: subbedByte=8'h5a;
		   8'h47: subbedByte=8'ha0;
		   8'h48: subbedByte=8'h52;
		   8'h49: subbedByte=8'h3b;
		   8'h4a: subbedByte=8'hd6;
		   8'h4b: subbedByte=8'hb3;
		   8'h4c: subbedByte=8'h29;
		   8'h4d: subbedByte=8'he3;
		   8'h4e: subbedByte=8'h2f;
		   8'h4f: subbedByte=8'h84;
		   8'h50: subbedByte=8'h53;
		   8'h51: subbedByte=8'hd1;
		   8'h52: subbedByte=8'h00;
		   8'h53: subbedByte=8'hed;
		   8'h54: subbedByte=8'h20;
		   8'h55: subbedByte=8'hfc;
		   8'h56: subbedByte=8'hb1;
		   8'h57: subbedByte=8'h5b;
		   8'h58: subbedByte=8'h6a;
		   8'h59: subbedByte=8'hcb;
		   8'h5a: subbedByte=8'hbe;
		   8'h5b: subbedByte=8'h39;
		   8'h5c: subbedByte=8'h4a;
		   8'h5d: subbedByte=8'h4c;
		   8'h5e: subbedByte=8'h58;
		   8'h5f: subbedByte=8'hcf;
		   8'h60: subbedByte=8'hd0;
		   8'h61: subbedByte=8'hef;
		   8'h62: subbedByte=8'haa;
		   8'h63: subbedByte=8'hfb;
		   8'h64: subbedByte=8'h43;
		   8'h65: subbedByte=8'h4d;
		   8'h66: subbedByte=8'h33;
		   8'h67: subbedByte=8'h85;
		   8'h68: subbedByte=8'h45;
		   8'h69: subbedByte=8'hf9;
		   8'h6a: subbedByte=8'h02;
		   8'h6b: subbedByte=8'h7f;
		   8'h6c: subbedByte=8'h50;
		   8'h6d: subbedByte=8'h3c;
		   8'h6e: subbedByte=8'h9f;
		   8'h6f: subbedByte=8'ha8;
		   8'h70: subbedByte=8'h51;
		   8'h71: subbedByte=8'ha3;
		   8'h72: subbedByte=8'h40;
		   8'h73: subbedByte=8'h8f;
		   8'h74: subbedByte=8'h92;
		   8'h75: subbedByte=8'h9d;
		   8'h76: subbedByte=8'h38;
		   8'h77: subbedByte=8'hf5;
		   8'h78: subbedByte=8'hbc;
		   8'h79: subbedByte=8'hb6;
		   8'h7a: subbedByte=8'hda;
		   8'h7b: subbedByte=8'h21;
		   8'h7c: subbedByte=8'h10;
		   8'h7d: subbedByte=8'hff;
		   8'h7e: subbedByte=8'hf3;
		   8'h7f: subbedByte=8'hd2;
		   8'h80: subbedByte=8'hcd;
		   8'h81: subbedByte=8'h0c;
		   8'h82: subbedByte=8'h13;
		   8'h83: subbedByte=8'hec;
		   8'h84: subbedByte=8'h5f;
		   8'h85: subbedByte=8'h97;
		   8'h86: subbedByte=8'h44;
		   8'h87: subbedByte=8'h17;
		   8'h88: subbedByte=8'hc4;
		   8'h89: subbedByte=8'ha7;
		   8'h8a: subbedByte=8'h7e;
		   8'h8b: subbedByte=8'h3d;
		   8'h8c: subbedByte=8'h64;
		   8'h8d: subbedByte=8'h5d;
		   8'h8e: subbedByte=8'h19;
		   8'h8f: subbedByte=8'h73;
		   8'h90: subbedByte=8'h60;
		   8'h91: subbedByte=8'h81;
		   8'h92: subbedByte=8'h4f;
		   8'h93: subbedByte=8'hdc;
		   8'h94: subbedByte=8'h22;
		   8'h95: subbedByte=8'h2a;
		   8'h96: subbedByte=8'h90;
		   8'h97: subbedByte=8'h88;
		   8'h98: subbedByte=8'h46;
		   8'h99: subbedByte=8'hee;
		   8'h9a: subbedByte=8'hb8;
		   8'h9b: subbedByte=8'h14;
		   8'h9c: subbedByte=8'hde;
		   8'h9d: subbedByte=8'h5e;
		   8'h9e: subbedByte=8'h0b;
		   8'h9f: subbedByte=8'hdb;
		   8'ha0: subbedByte=8'he0;
		   8'ha1: subbedByte=8'h32;
		   8'ha2: subbedByte=8'h3a;
		   8'ha3: subbedByte=8'h0a;
		   8'ha4: subbedByte=8'h49;
		   8'ha5: subbedByte=8'h06;
		   8'ha6: subbedByte=8'h24;
		   8'ha7: subbedByte=8'h5c;
		   8'ha8: subbedByte=8'hc2;
		   8'ha9: subbedByte=8'hd3;
		   8'haa: subbedByte=8'hac;
		   8'hab: subbedByte=8'h62;
		   8'hac: subbedByte=8'h91;
		   8'had: subbedByte=8'h95;
		   8'hae: subbedByte=8'he4;
		   8'haf: subbedByte=8'h79;
		   8'hb0: subbedByte=8'he7;
		   8'hb1: subbedByte=8'hc8;
		   8'hb2: subbedByte=8'h37;
		   8'hb3: subbedByte=8'h6d;
		   8'hb4: subbedByte=8'h8d;
		   8'hb5: subbedByte=8'hd5;
		   8'hb6: subbedByte=8'h4e;
		   8'hb7: subbedByte=8'ha9;
		   8'hb8: subbedByte=8'h6c;
		   8'hb9: subbedByte=8'h56;
		   8'hba: subbedByte=8'hf4;
		   8'hbb: subbedByte=8'hea;
		   8'hbc: subbedByte=8'h65;
		   8'hbd: subbedByte=8'h7a;
		   8'hbe: subbedByte=8'hae;
		   8'hbf: subbedByte=8'h08;
		   8'hc0: subbedByte=8'hba;
		   8'hc1: subbedByte=8'h78;
		   8'hc2: subbedByte=8'h25;
		   8'hc3: subbedByte=8'h2e;
		   8'hc4: subbedByte=8'h1c;
		   8'hc5: subbedByte=8'ha6;
		   8'hc6: subbedByte=8'hb4;
		   8'hc7: subbedByte=8'hc6;
		   8'hc8: subbedByte=8'he8;
		   8'hc9: subbedByte=8'hdd;
		   8'hca: subbedByte=8'h74;
		   8'hcb: subbedByte=8'h1f;
		   8'hcc: subbedByte=8'h4b;
		   8'hcd: subbedByte=8'hbd;
		   8'hce: subbedByte=8'h8b;
		   8'hcf: subbedByte=8'h8a;
		   8'hd0: subbedByte=8'h70;
		   8'hd1: subbedByte=8'h3e;
		   8'hd2: subbedByte=8'hb5;
		   8'hd3: subbedByte=8'h66;
		   8'hd4: subbedByte=8'h48;
		   8'hd5: subbedByte=8'h03;
		   8'hd6: subbedByte=8'hf6;
		   8'hd7: subbedByte=8'h0e;
		   8'hd8: subbedByte=8'h61;
		   8'hd9: subbedByte=8'h35;
		   8'hda: subbedByte=8'h57;
		   8'hdb: subbedByte=8'hb9;
		   8'hdc: subbedByte=8'h86;
		   8'hdd: subbedByte=8'hc1;
		   8'hde: subbedByte=8'h1d;
		   8'hdf: subbedByte=8'h9e;
		   8'he0: subbedByte=8'he1;
		   8'he1: subbedByte=8'hf8;
		   8'he2: subbedByte=8'h98;
		   8'he3: subbedByte=8'h11;
		   8'he4: subbedByte=8'h69;
		   8'he5: subbedByte=8'hd9;
		   8'he6: subbedByte=8'h8e;
		   8'he7: subbedByte=8'h94;
		   8'he8: subbedByte=8'h9b;
		   8'he9: subbedByte=8'h1e;
		   8'hea: subbedByte=8'h87;
		   8'heb: subbedByte=8'he9;
		   8'hec: subbedByte=8'hce;
		   8'hed: subbedByte=8'h55;
		   8'hee: subbedByte=8'h28;
		   8'hef: subbedByte=8'hdf;
		   8'hf0: subbedByte=8'h8c;
		   8'hf1: subbedByte=8'ha1;
		   8'hf2: subbedByte=8'h89;
		   8'hf3: subbedByte=8'h0d;
		   8'hf4: subbedByte=8'hbf;
		   8'hf5: subbedByte=8'he6;
		   8'hf6: subbedByte=8'h42;
		   8'hf7: subbedByte=8'h68;
		   8'hf8: subbedByte=8'h41;
		   8'hf9: subbedByte=8'h99;
		   8'hfa: subbedByte=8'h2d;
		   8'hfb: subbedByte=8'h0f;
		   8'hfc: subbedByte=8'hb0;
		   8'hfd: subbedByte=8'h54;
		   8'hfe: subbedByte=8'hbb;
		   8'hff: subbedByte=8'h16;
		endcase
    end
endmodule

