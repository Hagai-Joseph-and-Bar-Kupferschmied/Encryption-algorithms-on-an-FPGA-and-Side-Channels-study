module VarTxt_input_AES #(
					CYPHER_SIZE = 128
				)
				(
					input clk,
					input ena,
					input reset,
					output reg [127:0] plainText,
					output reg [CYPHER_SIZE-1:0] cypher_key
				);
	

	reg [6:0] idx; 
	
	always @(posedge clk or posedge reset)
	begin
		if (reset) begin
			plainText <= 0;
			cypher_key <= 0;
			idx <= 0;
		end
		else if (ena) begin
			plainText <= GenText(idx);
			cypher_key <= GenCKey(idx);
			idx <= idx + 1;
		end
	end


	function[127:0] GenText;
	input [6:0] idx;
	begin
	 case(idx)
		// VarTxt Test
		0: GenText = 128'h80000000000000000000000000000000;
		1: GenText = 128'hc0000000000000000000000000000000;
		2: GenText = 128'he0000000000000000000000000000000;
		3: GenText = 128'hf0000000000000000000000000000000;
		4: GenText = 128'hf8000000000000000000000000000000;
		5: GenText = 128'hfc000000000000000000000000000000;
		6: GenText = 128'hfe000000000000000000000000000000;
		7: GenText = 128'hff000000000000000000000000000000;
		8: GenText = 128'hff800000000000000000000000000000;
		9: GenText = 128'hffc00000000000000000000000000000;
		10: GenText = 128'hffe00000000000000000000000000000;
		11: GenText = 128'hfff00000000000000000000000000000;
		12: GenText = 128'hfff80000000000000000000000000000;
		13: GenText = 128'hfffc0000000000000000000000000000;
		14: GenText = 128'hfffe0000000000000000000000000000;
		15: GenText = 128'hffff0000000000000000000000000000;
		16: GenText = 128'hffff8000000000000000000000000000;
		17: GenText = 128'hffffc000000000000000000000000000;
		18: GenText = 128'hffffe000000000000000000000000000;
		19: GenText = 128'hfffff000000000000000000000000000;
		20: GenText = 128'hfffff800000000000000000000000000;
		21: GenText = 128'hfffffc00000000000000000000000000;
		22: GenText = 128'hfffffe00000000000000000000000000;
		23: GenText = 128'hffffff00000000000000000000000000;
		24: GenText = 128'hffffff80000000000000000000000000;
		25: GenText = 128'hffffffc0000000000000000000000000;
		26: GenText = 128'hffffffe0000000000000000000000000;
		27: GenText = 128'hfffffff0000000000000000000000000;
		28: GenText = 128'hfffffff8000000000000000000000000;
		29: GenText = 128'hfffffffc000000000000000000000000;
		30: GenText = 128'hfffffffe000000000000000000000000;
		31: GenText = 128'hffffffff000000000000000000000000;
		32: GenText = 128'hffffffff800000000000000000000000;
		33: GenText = 128'hffffffffc00000000000000000000000;
		34: GenText = 128'hffffffffe00000000000000000000000;
		35: GenText = 128'hfffffffff00000000000000000000000;
		36: GenText = 128'hfffffffff80000000000000000000000;
		37: GenText = 128'hfffffffffc0000000000000000000000;
		38: GenText = 128'hfffffffffe0000000000000000000000;
		39: GenText = 128'hffffffffff0000000000000000000000;
		40: GenText = 128'hffffffffff8000000000000000000000;
		41: GenText = 128'hffffffffffc000000000000000000000;
		42: GenText = 128'hffffffffffe000000000000000000000;
		43: GenText = 128'hfffffffffff000000000000000000000;
		44: GenText = 128'hfffffffffff800000000000000000000;
		45: GenText = 128'hfffffffffffc00000000000000000000;
		46: GenText = 128'hfffffffffffe00000000000000000000;
		47: GenText = 128'hffffffffffff00000000000000000000;
		48: GenText = 128'hffffffffffff80000000000000000000;
		49: GenText = 128'hffffffffffffc0000000000000000000;
		50: GenText = 128'hffffffffffffe0000000000000000000;
		51: GenText = 128'hfffffffffffff0000000000000000000;
		52: GenText = 128'hfffffffffffff8000000000000000000;
		53: GenText = 128'hfffffffffffffc000000000000000000;
		54: GenText = 128'hfffffffffffffe000000000000000000;
		55: GenText = 128'hffffffffffffff000000000000000000;
		56: GenText = 128'hffffffffffffff800000000000000000;
		57: GenText = 128'hffffffffffffffc00000000000000000;
		58: GenText = 128'hffffffffffffffe00000000000000000;
		59: GenText = 128'hfffffffffffffff00000000000000000;
		60: GenText = 128'hfffffffffffffff80000000000000000;
		61: GenText = 128'hfffffffffffffffc0000000000000000;
		62: GenText = 128'hfffffffffffffffe0000000000000000;
		63: GenText = 128'hffffffffffffffff0000000000000000;
		64: GenText = 128'hffffffffffffffff8000000000000000;
		65: GenText = 128'hffffffffffffffffc000000000000000;
		66: GenText = 128'hffffffffffffffffe000000000000000;
		67: GenText = 128'hfffffffffffffffff000000000000000;
		68: GenText = 128'hfffffffffffffffff800000000000000;
		69: GenText = 128'hfffffffffffffffffc00000000000000;
		70: GenText = 128'hfffffffffffffffffe00000000000000;
		71: GenText = 128'hffffffffffffffffff00000000000000;
		72: GenText = 128'hffffffffffffffffff80000000000000;
		73: GenText = 128'hffffffffffffffffffc0000000000000;
		74: GenText = 128'hffffffffffffffffffe0000000000000;
		75: GenText = 128'hfffffffffffffffffff0000000000000;
		76: GenText = 128'hfffffffffffffffffff8000000000000;
		77: GenText = 128'hfffffffffffffffffffc000000000000;
		78: GenText = 128'hfffffffffffffffffffe000000000000;
		79: GenText = 128'hffffffffffffffffffff000000000000;
		80: GenText = 128'hffffffffffffffffffff800000000000;
		81: GenText = 128'hffffffffffffffffffffc00000000000;
		82: GenText = 128'hffffffffffffffffffffe00000000000;
		83: GenText = 128'hfffffffffffffffffffff00000000000;
		84: GenText = 128'hfffffffffffffffffffff80000000000;
		85: GenText = 128'hfffffffffffffffffffffc0000000000;
		86: GenText = 128'hfffffffffffffffffffffe0000000000;
		87: GenText = 128'hffffffffffffffffffffff0000000000;
		88: GenText = 128'hffffffffffffffffffffff8000000000;
		89: GenText = 128'hffffffffffffffffffffffc000000000;
		90: GenText = 128'hffffffffffffffffffffffe000000000;
		91: GenText = 128'hfffffffffffffffffffffff000000000;
		92: GenText = 128'hfffffffffffffffffffffff800000000;
		93: GenText = 128'hfffffffffffffffffffffffc00000000;
		94: GenText = 128'hfffffffffffffffffffffffe00000000;
		95: GenText = 128'hffffffffffffffffffffffff00000000;
		96: GenText = 128'hffffffffffffffffffffffff80000000;
		97: GenText = 128'hffffffffffffffffffffffffc0000000;
		98: GenText = 128'hffffffffffffffffffffffffe0000000;
		99: GenText = 128'hfffffffffffffffffffffffff0000000;
		100: GenText = 128'hfffffffffffffffffffffffff8000000;
		101: GenText = 128'hfffffffffffffffffffffffffc000000;
		102: GenText = 128'hfffffffffffffffffffffffffe000000;
		103: GenText = 128'hffffffffffffffffffffffffff000000;
		104: GenText = 128'hffffffffffffffffffffffffff800000;
		105: GenText = 128'hffffffffffffffffffffffffffc00000;
		106: GenText = 128'hffffffffffffffffffffffffffe00000;
		107: GenText = 128'hfffffffffffffffffffffffffff00000;
		108: GenText = 128'hfffffffffffffffffffffffffff80000;
		109: GenText = 128'hfffffffffffffffffffffffffffc0000;
		110: GenText = 128'hfffffffffffffffffffffffffffe0000;
		111: GenText = 128'hffffffffffffffffffffffffffff0000;
		112: GenText = 128'hffffffffffffffffffffffffffff8000;
		113: GenText = 128'hffffffffffffffffffffffffffffc000;
		114: GenText = 128'hffffffffffffffffffffffffffffe000;
		115: GenText = 128'hfffffffffffffffffffffffffffff000;
		116: GenText = 128'hfffffffffffffffffffffffffffff800;
		117: GenText = 128'hfffffffffffffffffffffffffffffc00;
		118: GenText = 128'hfffffffffffffffffffffffffffffe00;
		119: GenText = 128'hffffffffffffffffffffffffffffff00;
		120: GenText = 128'hffffffffffffffffffffffffffffff80;
		121: GenText = 128'hffffffffffffffffffffffffffffffc0;
		122: GenText = 128'hffffffffffffffffffffffffffffffe0;
		123: GenText = 128'hfffffffffffffffffffffffffffffff0;
		124: GenText = 128'hfffffffffffffffffffffffffffffff8;
		125: GenText = 128'hfffffffffffffffffffffffffffffffc;
		126: GenText = 128'hfffffffffffffffffffffffffffffffe;
		127: GenText = 128'hffffffffffffffffffffffffffffffff;
		default: GenText = 0;
	  endcase
	  end
	endfunction
	
	function[CYPHER_SIZE-1:0] GenCKey;
	input [6:0] idx; 
	begin
	 case(idx)
		// VarTxt Test
		0: GenCKey = 128'h00000000000000000000000000000000;
		1: GenCKey = 128'h00000000000000000000000000000000;
		2: GenCKey = 128'h00000000000000000000000000000000;
		3: GenCKey = 128'h00000000000000000000000000000000;
		4: GenCKey = 128'h00000000000000000000000000000000;
		5: GenCKey = 128'h00000000000000000000000000000000;
		6: GenCKey = 128'h00000000000000000000000000000000;
		7: GenCKey = 128'h00000000000000000000000000000000;
		8: GenCKey = 128'h00000000000000000000000000000000;
		9: GenCKey = 128'h00000000000000000000000000000000;
		10: GenCKey = 128'h00000000000000000000000000000000;
		11: GenCKey = 128'h00000000000000000000000000000000;
		12: GenCKey = 128'h00000000000000000000000000000000;
		13: GenCKey = 128'h00000000000000000000000000000000;
		14: GenCKey = 128'h00000000000000000000000000000000;
		15: GenCKey = 128'h00000000000000000000000000000000;
		16: GenCKey = 128'h00000000000000000000000000000000;
		17: GenCKey = 128'h00000000000000000000000000000000;
		18: GenCKey = 128'h00000000000000000000000000000000;
		19: GenCKey = 128'h00000000000000000000000000000000;
		20: GenCKey = 128'h00000000000000000000000000000000;
		21: GenCKey = 128'h00000000000000000000000000000000;
		22: GenCKey = 128'h00000000000000000000000000000000;
		23: GenCKey = 128'h00000000000000000000000000000000;
		24: GenCKey = 128'h00000000000000000000000000000000;
		25: GenCKey = 128'h00000000000000000000000000000000;
		26: GenCKey = 128'h00000000000000000000000000000000;
		27: GenCKey = 128'h00000000000000000000000000000000;
		28: GenCKey = 128'h00000000000000000000000000000000;
		29: GenCKey = 128'h00000000000000000000000000000000;
		30: GenCKey = 128'h00000000000000000000000000000000;
		31: GenCKey = 128'h00000000000000000000000000000000;
		32: GenCKey = 128'h00000000000000000000000000000000;
		33: GenCKey = 128'h00000000000000000000000000000000;
		34: GenCKey = 128'h00000000000000000000000000000000;
		35: GenCKey = 128'h00000000000000000000000000000000;
		36: GenCKey = 128'h00000000000000000000000000000000;
		37: GenCKey = 128'h00000000000000000000000000000000;
		38: GenCKey = 128'h00000000000000000000000000000000;
		39: GenCKey = 128'h00000000000000000000000000000000;
		40: GenCKey = 128'h00000000000000000000000000000000;
		41: GenCKey = 128'h00000000000000000000000000000000;
		42: GenCKey = 128'h00000000000000000000000000000000;
		43: GenCKey = 128'h00000000000000000000000000000000;
		44: GenCKey = 128'h00000000000000000000000000000000;
		45: GenCKey = 128'h00000000000000000000000000000000;
		46: GenCKey = 128'h00000000000000000000000000000000;
		47: GenCKey = 128'h00000000000000000000000000000000;
		48: GenCKey = 128'h00000000000000000000000000000000;
		49: GenCKey = 128'h00000000000000000000000000000000;
		50: GenCKey = 128'h00000000000000000000000000000000;
		51: GenCKey = 128'h00000000000000000000000000000000;
		52: GenCKey = 128'h00000000000000000000000000000000;
		53: GenCKey = 128'h00000000000000000000000000000000;
		54: GenCKey = 128'h00000000000000000000000000000000;
		55: GenCKey = 128'h00000000000000000000000000000000;
		56: GenCKey = 128'h00000000000000000000000000000000;
		57: GenCKey = 128'h00000000000000000000000000000000;
		58: GenCKey = 128'h00000000000000000000000000000000;
		59: GenCKey = 128'h00000000000000000000000000000000;
		60: GenCKey = 128'h00000000000000000000000000000000;
		61: GenCKey = 128'h00000000000000000000000000000000;
		62: GenCKey = 128'h00000000000000000000000000000000;
		63: GenCKey = 128'h00000000000000000000000000000000;
		64: GenCKey = 128'h00000000000000000000000000000000;
		65: GenCKey = 128'h00000000000000000000000000000000;
		66: GenCKey = 128'h00000000000000000000000000000000;
		67: GenCKey = 128'h00000000000000000000000000000000;
		68: GenCKey = 128'h00000000000000000000000000000000;
		69: GenCKey = 128'h00000000000000000000000000000000;
		70: GenCKey = 128'h00000000000000000000000000000000;
		71: GenCKey = 128'h00000000000000000000000000000000;
		72: GenCKey = 128'h00000000000000000000000000000000;
		73: GenCKey = 128'h00000000000000000000000000000000;
		74: GenCKey = 128'h00000000000000000000000000000000;
		75: GenCKey = 128'h00000000000000000000000000000000;
		76: GenCKey = 128'h00000000000000000000000000000000;
		77: GenCKey = 128'h00000000000000000000000000000000;
		78: GenCKey = 128'h00000000000000000000000000000000;
		79: GenCKey = 128'h00000000000000000000000000000000;
		80: GenCKey = 128'h00000000000000000000000000000000;
		81: GenCKey = 128'h00000000000000000000000000000000;
		82: GenCKey = 128'h00000000000000000000000000000000;
		83: GenCKey = 128'h00000000000000000000000000000000;
		84: GenCKey = 128'h00000000000000000000000000000000;
		85: GenCKey = 128'h00000000000000000000000000000000;
		86: GenCKey = 128'h00000000000000000000000000000000;
		87: GenCKey = 128'h00000000000000000000000000000000;
		88: GenCKey = 128'h00000000000000000000000000000000;
		89: GenCKey = 128'h00000000000000000000000000000000;
		90: GenCKey = 128'h00000000000000000000000000000000;
		91: GenCKey = 128'h00000000000000000000000000000000;
		92: GenCKey = 128'h00000000000000000000000000000000;
		93: GenCKey = 128'h00000000000000000000000000000000;
		94: GenCKey = 128'h00000000000000000000000000000000;
		95: GenCKey = 128'h00000000000000000000000000000000;
		96: GenCKey = 128'h00000000000000000000000000000000;
		97: GenCKey = 128'h00000000000000000000000000000000;
		98: GenCKey = 128'h00000000000000000000000000000000;
		99: GenCKey = 128'h00000000000000000000000000000000;
		100: GenCKey = 128'h00000000000000000000000000000000;
		101: GenCKey = 128'h00000000000000000000000000000000;
		102: GenCKey = 128'h00000000000000000000000000000000;
		103: GenCKey = 128'h00000000000000000000000000000000;
		104: GenCKey = 128'h00000000000000000000000000000000;
		105: GenCKey = 128'h00000000000000000000000000000000;
		106: GenCKey = 128'h00000000000000000000000000000000;
		107: GenCKey = 128'h00000000000000000000000000000000;
		108: GenCKey = 128'h00000000000000000000000000000000;
		109: GenCKey = 128'h00000000000000000000000000000000;
		110: GenCKey = 128'h00000000000000000000000000000000;
		111: GenCKey = 128'h00000000000000000000000000000000;
		112: GenCKey = 128'h00000000000000000000000000000000;
		113: GenCKey = 128'h00000000000000000000000000000000;
		114: GenCKey = 128'h00000000000000000000000000000000;
		115: GenCKey = 128'h00000000000000000000000000000000;
		116: GenCKey = 128'h00000000000000000000000000000000;
		117: GenCKey = 128'h00000000000000000000000000000000;
		118: GenCKey = 128'h00000000000000000000000000000000;
		119: GenCKey = 128'h00000000000000000000000000000000;
		120: GenCKey = 128'h00000000000000000000000000000000;
		121: GenCKey = 128'h00000000000000000000000000000000;
		122: GenCKey = 128'h00000000000000000000000000000000;
		123: GenCKey = 128'h00000000000000000000000000000000;
		124: GenCKey = 128'h00000000000000000000000000000000;
		125: GenCKey = 128'h00000000000000000000000000000000;
		126: GenCKey = 128'h00000000000000000000000000000000;
		127: GenCKey = 128'h00000000000000000000000000000000;
		default: GenCKey = 0;
	  endcase
	  end
	endfunction
	
endmodule